CONFIGURATION ControlUnit_Behavior_config OF ControlUnit IS
   FOR Behavior
   END FOR;
END ControlUnit_Behavior_config;