--
-- VHDL Architecture ADD_SingleCycle_lib.ent.arch
--
-- Created:
--          by - jwarchal.UNKNOWN (GURREN)
--          at - 12:13:46 02/ 1/2013
--
-- using Mentor Graphics HDL Designer(TM) 2012.1 (Build 6)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY ent IS
END ENTITY ent;

--
ARCHITECTURE arch OF ent IS
BEGIN
END ARCHITECTURE arch;

