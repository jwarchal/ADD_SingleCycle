CONFIGURATION mux2to1_mux2to1arch_config OF mux2to1 IS
   FOR mux2to1arch
   END FOR;
END mux2to1_mux2to1arch_config;