CONFIGURATION Extendblock_Extendblockarch_config OF Extendblock IS
   FOR Extendblockarch
   END FOR;
END Extendblock_Extendblockarch_config;