CONFIGURATION PC_PCarch_config OF PC IS
   FOR PCarch
   END FOR;
END PC_PCarch_config;