CONFIGURATION alu_aluarch_config OF alu IS
   FOR aluarch
   END FOR;
END alu_aluarch_config;