CONFIGURATION RegisterFile_Behavior_config OF RegisterFile IS
   FOR Behavior
   END FOR;
END RegisterFile_Behavior_config;