--
-- VHDL Architecture ADD_SingleCycle_lib.Increment.Incrementarch
--
-- Created:
--          by - Vincent.UNKNOWN (VINCENT-LAPTOP)
--          at - 15:42:19 02/ 5/2013
--
-- using Mentor Graphics HDL Designer(TM) 2012.1 (Build 6)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY Increment IS
  PORT(a: IN std_logic_vector(15 DOWNTO 0);
    b: OUT std_logic_vector(15 DOWNTO 0));
END ENTITY Increment;

--
ARCHITECTURE Incrementarch OF Increment IS
  BEGIN
  PROCESS(a)
  CONSTANT one: unsigned(15 DOWNTO 0):= "0000000000000001";
  VARIABLE locala: unsigned(15 DOWNTO 0);
  VARIABLE localb: unsigned(15 DOWNTO 0);
  BEGIN
    locala:= unsigned(a(15 DOWNTO 0));
    localb:= (locala + one);
    b <= std_logic_vector(localb);
END PROCESS;
END ARCHITECTURE Incrementarch;

