CONFIGURATION mux4to1_mux4to1arch_config OF mux4to1 IS
   FOR mux4to1arch
   END FOR;
END mux4to1_mux4to1arch_config;