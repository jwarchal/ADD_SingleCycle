CONFIGURATION Increment_Incrementarch_config OF Increment IS
   FOR Incrementarch
   END FOR;
END Increment_Incrementarch_config;